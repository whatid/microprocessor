library verilog;
use verilog.vl_types.all;
entity instructionMem_sv_unit is
end instructionMem_sv_unit;
