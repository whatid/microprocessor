library verilog;
use verilog.vl_types.all;
entity ControlROM_sv_unit is
end ControlROM_sv_unit;
