library verilog;
use verilog.vl_types.all;
entity mux5_sv_unit is
end mux5_sv_unit;
