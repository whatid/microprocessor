library verilog;
use verilog.vl_types.all;
entity branch_logic_sv_unit is
end branch_logic_sv_unit;
