library verilog;
use verilog.vl_types.all;
entity pc_array_sv_unit is
end pc_array_sv_unit;
