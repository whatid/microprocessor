library verilog;
use verilog.vl_types.all;
entity mp3_mod_sv_unit is
end mp3_mod_sv_unit;
