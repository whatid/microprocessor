library verilog;
use verilog.vl_types.all;
entity lru_array_sv_unit is
end lru_array_sv_unit;
