library verilog;
use verilog.vl_types.all;
entity zextshift_sv_unit is
end zextshift_sv_unit;
