library verilog;
use verilog.vl_types.all;
entity L2_tagmux_sv_unit is
end L2_tagmux_sv_unit;
