library verilog;
use verilog.vl_types.all;
entity L2_Cache_sv_unit is
end L2_Cache_sv_unit;
