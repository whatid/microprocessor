library verilog;
use verilog.vl_types.all;
entity data_sv_unit is
end data_sv_unit;
