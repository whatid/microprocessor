library verilog;
use verilog.vl_types.all;
entity instructionWB_sv_unit is
end instructionWB_sv_unit;
