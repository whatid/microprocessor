library verilog;
use verilog.vl_types.all;
entity datamux_sv_unit is
end datamux_sv_unit;
