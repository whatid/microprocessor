library verilog;
use verilog.vl_types.all;
entity InstructionExecute_sv_unit is
end InstructionExecute_sv_unit;
