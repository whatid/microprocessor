library verilog;
use verilog.vl_types.all;
entity InstructionDecode_sv_unit is
end InstructionDecode_sv_unit;
