library verilog;
use verilog.vl_types.all;
entity hazard_detection_sv_unit is
end hazard_detection_sv_unit;
