library verilog;
use verilog.vl_types.all;
entity L2_cache_control_sv_unit is
end L2_cache_control_sv_unit;
