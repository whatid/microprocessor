library verilog;
use verilog.vl_types.all;
entity L2_cache_datapath is
    port(
        clk             : in     vl_logic;
        write_back      : in     vl_logic;
        write1          : in     vl_logic;
        write2          : in     vl_logic;
        write3          : in     vl_logic;
        write4          : in     vl_logic;
        way1            : in     vl_logic;
        way2            : in     vl_logic;
        way3            : in     vl_logic;
        way4            : in     vl_logic;
        load_dbit1      : in     vl_logic;
        load_dbit2      : in     vl_logic;
        load_dbit3      : in     vl_logic;
        load_dbit4      : in     vl_logic;
        set_dbit        : in     vl_logic;
        set_vbit        : in     vl_logic;
        load_vbit1      : in     vl_logic;
        load_vbit2      : in     vl_logic;
        load_vbit3      : in     vl_logic;
        load_vbit4      : in     vl_logic;
        load_data1      : in     vl_logic;
        load_data2      : in     vl_logic;
        load_data3      : in     vl_logic;
        load_data4      : in     vl_logic;
        load_tag1       : in     vl_logic;
        load_tag2       : in     vl_logic;
        load_tag3       : in     vl_logic;
        load_tag4       : in     vl_logic;
        data_sel        : in     vl_logic_vector(1 downto 0);
        phys_sel        : in     vl_logic_vector(1 downto 0);
        lru_out         : out    vl_logic_vector(1 downto 0);
        dirty_out1      : out    vl_logic;
        dirty_out2      : out    vl_logic;
        dirty_out3      : out    vl_logic;
        dirty_out4      : out    vl_logic;
        access1         : out    vl_logic;
        access2         : out    vl_logic;
        access3         : out    vl_logic;
        access4         : out    vl_logic;
        hit             : out    vl_logic;
        mem_address     : in     vl_logic_vector(15 downto 0);
        pmem_rdata      : in     vl_logic_vector(127 downto 0);
        mem_wdata       : in     vl_logic_vector(127 downto 0);
        pmem_wdata      : out    vl_logic_vector(127 downto 0);
        mem_rdata       : out    vl_logic_vector(127 downto 0);
        pmem_address    : out    vl_logic_vector(15 downto 0)
    );
end L2_cache_datapath;
