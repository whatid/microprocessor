library verilog;
use verilog.vl_types.all;
entity adder_sv_unit is
end adder_sv_unit;
