library verilog;
use verilog.vl_types.all;
entity tag_comparator_sv_unit is
end tag_comparator_sv_unit;
