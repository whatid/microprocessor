library verilog;
use verilog.vl_types.all;
entity instr_array_sv_unit is
end instr_array_sv_unit;
