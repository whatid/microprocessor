library verilog;
use verilog.vl_types.all;
entity address_parser_sv_unit is
end address_parser_sv_unit;
