library verilog;
use verilog.vl_types.all;
entity btb_sv_unit is
end btb_sv_unit;
