library verilog;
use verilog.vl_types.all;
entity tagmux_sv_unit is
end tagmux_sv_unit;
