library verilog;
use verilog.vl_types.all;
entity mux3_sv_unit is
end mux3_sv_unit;
