library verilog;
use verilog.vl_types.all;
entity InstructionFetch_sv_unit is
end InstructionFetch_sv_unit;
