library verilog;
use verilog.vl_types.all;
entity L2_cache_control is
    port(
        clk             : in     vl_logic;
        lru_out         : in     vl_logic_vector(1 downto 0);
        dirty_out1      : in     vl_logic;
        dirty_out2      : in     vl_logic;
        dirty_out3      : in     vl_logic;
        dirty_out4      : in     vl_logic;
        access1         : in     vl_logic;
        access2         : in     vl_logic;
        access3         : in     vl_logic;
        access4         : in     vl_logic;
        way1            : out    vl_logic;
        way2            : out    vl_logic;
        way3            : out    vl_logic;
        way4            : out    vl_logic;
        hit             : in     vl_logic;
        write1          : out    vl_logic;
        write2          : out    vl_logic;
        write3          : out    vl_logic;
        write4          : out    vl_logic;
        load_dbit1      : out    vl_logic;
        load_dbit2      : out    vl_logic;
        load_dbit3      : out    vl_logic;
        load_dbit4      : out    vl_logic;
        set_dbit        : out    vl_logic;
        set_vbit        : out    vl_logic;
        load_vbit1      : out    vl_logic;
        load_vbit2      : out    vl_logic;
        load_vbit3      : out    vl_logic;
        load_vbit4      : out    vl_logic;
        load_data1      : out    vl_logic;
        load_data2      : out    vl_logic;
        load_data3      : out    vl_logic;
        load_data4      : out    vl_logic;
        load_tag1       : out    vl_logic;
        load_tag2       : out    vl_logic;
        load_tag3       : out    vl_logic;
        load_tag4       : out    vl_logic;
        data_sel        : out    vl_logic_vector(1 downto 0);
        write_back      : out    vl_logic;
        phys_sel        : out    vl_logic_vector(1 downto 0);
        mem_read        : in     vl_logic;
        mem_write       : in     vl_logic;
        pmem_resp       : in     vl_logic;
        pmem_read       : out    vl_logic;
        pmem_write      : out    vl_logic;
        mem_resp        : out    vl_logic
    );
end L2_cache_control;
