library verilog;
use verilog.vl_types.all;
entity decoder_sv_unit is
end decoder_sv_unit;
