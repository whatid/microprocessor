library verilog;
use verilog.vl_types.all;
entity mp3_datapath_sv_unit is
end mp3_datapath_sv_unit;
