module andgate
(
	input logic a,
	input logic b,
	output c
);

assign c = a && b; 

endmodule : andgate 
