library verilog;
use verilog.vl_types.all;
entity mux4_sv_unit is
end mux4_sv_unit;
