library verilog;
use verilog.vl_types.all;
entity comparator_sv_unit is
end comparator_sv_unit;
