library verilog;
use verilog.vl_types.all;
entity L2_address_parser_sv_unit is
end L2_address_parser_sv_unit;
