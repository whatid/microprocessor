library verilog;
use verilog.vl_types.all;
entity counter_sv_unit is
end counter_sv_unit;
