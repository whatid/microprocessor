library verilog;
use verilog.vl_types.all;
entity mp3 is
end mp3;
