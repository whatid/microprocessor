library verilog;
use verilog.vl_types.all;
entity trim_byte_sv_unit is
end trim_byte_sv_unit;
