library verilog;
use verilog.vl_types.all;
entity arbiter_datapath_sv_unit is
end arbiter_datapath_sv_unit;
