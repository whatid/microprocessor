library verilog;
use verilog.vl_types.all;
entity ID_Datapath_sv_unit is
end ID_Datapath_sv_unit;
